module FIR(x, y, clk, reset);



endmodule
